library ieee;
use ieee.std_logic_1164.all;

entity top is
    port (
        tram_wr_en : in  std_logic;
        reset      : in  std_logic;
        clk_48     : out std_logic;
        clk_tx     : out std_logic;
        dout       : out std_logic;
        enc_ena    : out std_logic
    );
end entity top;

architecture rtl of top is
    component tx_tb is
        generic (
            BITS      :     INTEGER := 10;           -- Number of bits being encoded
            mlength   :     INTEGER := 11            -- Number of bits in the length message (not including the sync)
        );
        port (
            wr_clk    : in  STD_LOGIC;
            reset     : in  STD_LOGIC;
            wr_en     : in  STD_LOGIC;
            tx_length : in  std_logic_vector(mlength - 1 downto 0);
            wr_ram    : out STD_LOGIC_VECTOR(BITS - 1 downto 0);
            wr_addr   : out STD_LOGIC_VECTOR(mlength - 1 downto 0);
            tx_ready  : out STD_LOGIC
        );
    end component tx_tb;

    component ram is
        generic (
            addr_width :     natural := 9;           -- 512x8
            data_width :     natural := 8
        );
        port (
            write_en   : in  std_logic;
            waddr      : in  std_logic_vector(addr_width - 1 downto 0);
            wclk       : in  std_logic;
            raddr      : in  std_logic_vector(addr_width - 1 downto 0);
            rclk       : in  std_logic;
            din        : in  std_logic_vector(data_width - 1 downto 0);
            dout       : out std_logic_vector(data_width - 1 downto 0)
        );
    end component ram;

    component manchester_encoder is
        generic (
            BITS         :     INTEGER := 10;        -- Number of bits being encoded
            mlength      :     INTEGER := 11         -- Number of bits in the length message (not including the sync)
        );
        port (
            clk          : in  STD_LOGIC;
            message      : in  STD_LOGIC_VECTOR(BITS - 1 downto 0);
            tx_length    : in  std_logic_vector(mlength - 1 downto 0);
            dout         : out STD_LOGIC;
            rd_addr      : out STD_LOGIC_VECTOR(mlength - 1 downto 0);
            message_sent : out STD_LOGIC;
            reset        : in  STD_LOGIC;
            ena_t        : in  STD_LOGIC
        );
    end component manchester_encoder;

    component clk_divider is
        generic (
            Freq_in :     INTEGER := 48000000;
            N       :     INTEGER := 10              -- speed divider, equates to the number of bits (BITS)
        );
        port (
            clk_in  : in  STD_LOGIC;
            reset   : in  STD_LOGIC;
            clk_out : out STD_LOGIC
        );
    end component clk_divider;


    component LT_controller is
        port (
            fsm_clk      : in  STD_LOGIC;
            rst          : in  STD_LOGIC;
            -- Indicators from other blocks to trigger states
            tx_ready     : in  STD_LOGIC;            -- indication from EC to start reading TX_RAM and transmit
            -- rx_received : IN STD_LOGIC; -- indication from the RX line that a light message is incoming
            -- host_align : IN STD_LOGIC;
            -- device_align : IN STD_LOGIC;
            -- Add error signals that suggest to go to idle state?
            -- rx_error : OUT STD_LOGIC;
            -- tx_error : OUT STD_LOGIC;
            -- host : IN STD_LOGIC;
            ena_t        : out std_logic;
            message_sent : in  std_logic
            -- rx_done : in std_logic;
            -- aligned : in std_logic
        );
    end component LT_controller;

    component SB_HFOSC is
        generic (
            CLKHF_DIV :     STRING := "0b00"
        );
        port (
            CLKHFEN   : in  STD_LOGIC;
            CLKHFPU   : in  STD_LOGIC;
            CLKHF     : out STD_LOGIC
        );
    end component SB_HFOSC;


    component SB_GB is
        port (
            USER_SIGNAL_TO_GLOBAL_BUFFER : in  std_logic;
            GLOBAL_BUFFER_OUTPUT         : out std_logic
        );
    end component SB_GB;

    signal tx_ready, tram_rd_en       : std_logic                     := '0';
    signal tram_in, tram_out          : std_logic_vector(11 downto 0);
    signal tx_clk                     : std_logic;
    signal tram_raddr_i, tram_waddr_i : std_logic_vector(10 downto 0);
    signal tx_length                  : std_logic_vector(10 downto 0) := "00001111111";
    signal ena_t                      : std_logic;
    signal message_sent               : std_logic                     := '0';
    signal enc_clk                    : std_logic;
    -- signal rx_received : std_logic := '0'; -- indication from the RX line that a light message is incoming
    -- signal host_align : std_logic := '0';
    -- signal device_align : std_logic := '0';
    -- 	-- Add error signals that suggest to go to idle state?
    -- signal rx_error : std_logic := '0';
    -- signal tx_error : std_logic := '0';
    -- signal host : std_logic := '0';
    -- signal rx_done : std_logic := '0';
    -- signal aligned : std_logic := '0';
    signal enc_clk_raw                : std_logic;
    signal enc_clk_glb                : std_logic;

begin
    tx_length <= "00000000111";

    ECin: component tx_tb
    generic map (
        BITS                         => 12,
        mlength                      => 11
    )
    port map (
        wr_clk                       => tx_clk,
        reset                        => reset,
        wr_en                        => tram_wr_en,
        tx_length                    => tx_length,
        wr_ram                       => tram_in,
        wr_addr                      => tram_waddr_i,
        tx_ready                     => tx_ready
    );

    ram_tx: component ram
    generic map (
        addr_width                   => 11,
        data_width                   => 12
    )
    port map (
        write_en                     => tram_wr_en,
        waddr                        => tram_waddr_i,
        wclk                         => tx_clk,
        raddr                        => tram_raddr_i,
        rclk                         => enc_clk_glb, -- **use global**
        din                          => tram_in,
        dout                         => tram_out
    );

    man_enc: component manchester_encoder
    generic map (
        BITS                         => 12,
        mlength                      => 11
    )
    port map (
        clk                          => enc_clk_glb, -- **use global**
        message                      => tram_out,
        tx_length                    => tx_length,
        dout                         => dout,
        rd_addr                      => tram_raddr_i,
        message_sent                 => message_sent,
        reset                        => reset,
        ena_t                        => ena_t
    );

    clk_4_tx: component clk_divider
    generic map (
        Freq_in                      => 48000000,
        N                            => 4
    )
    port map (
        clk_in                       => enc_clk_glb, -- **use global**
        reset                        => reset,
        clk_out                      => tx_clk
    );

    lt_fsm: component LT_controller
    port map (
        fsm_clk                      => enc_clk_glb, -- **use global**
        rst                          => reset,
        tx_ready                     => tx_ready,
        ena_t                        => ena_t,
        message_sent                 => message_sent
    );

    -- HFOSC -> raw clock
    u_osc: component SB_HFOSC
    generic map (
        CLKHF_DIV                    => "0b00"
    )
    port map (
        CLKHFEN                      => '1',
        CLKHFPU                      => '1',
        CLKHF                        => enc_clk_raw
    );

    -- >>> NEW: global buffer for 48 MHz domain
    u_clk48_gb: component SB_GB
    port map (
        USER_SIGNAL_TO_GLOBAL_BUFFER => enc_clk_raw,
        GLOBAL_BUFFER_OUTPUT         => enc_clk_glb
    );
    -- <<<

    -- Outputs
    clk_48    <= enc_clk_glb;                        -- expose the global’d clock
    clk_tx    <= tx_clk;
    enc_ena   <= ena_t;

end architecture rtl;
